`timescale 1ns / 1ps

module OR(
input I1,I2,
output O
    );
    
    assign O=I1||I2;
    
endmodule
