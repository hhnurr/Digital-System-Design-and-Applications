`timescale 1ns / 1ps

module NOT(

input I,
output O

    );
    
   assign O=~I;
endmodule
