`timescale 1ns / 1ps

module AND(
input I1,I2,
output O
    );
    
    assign O=I1&I2;
    
endmodule
